module top_module (
    input ring,
    input vibrate_mode,
    output ringer,       // Make sound
    output motor         // Vibrate
);
    assign ringer = ring ^ motor;
	assign motor = vibrate_mode & ring;
    

endmodule
