module top_module(output zero);
    /*atribuindo = <largura, base, valor>*/
    assign zero = 1'b0;

endmodule
