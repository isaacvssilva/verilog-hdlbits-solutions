module top_module(output one);
    /*atribuindo = <largura, base, valor>*/
    assign one = 1'b1;
endmodule
