module top_module(input in, output out);
    /*input in --wire--> output out */
	assign out = in;
endmodule
